// Multi-input AND gate
module red(input [3:0] i, output o);
  assign o = &i;
endmodule

