// high impedance state
module sourceZ(
  output out
);
  assign out = 1'bZ;

endmodule